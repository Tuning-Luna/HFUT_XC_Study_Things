// ============================================================================
// 指令存储器模块
// ============================================================================
// 功能：存储程序指令，根据地址读取指令
// 输入：addr - 指令地址（PC 值）
// 输出：instruction - 32 位指令
// 说明：本模块预装载了6条指令测试程序（add, sub, and, or, slt, addi）
// ============================================================================

`timescale 1ns/1ps

module instruction_memory(
    input wire [31:0] addr,          // 指令地址
    output wire [31:0] instruction   // 输出指令
);

    // 指令存储器（128 条指令）
    reg [31:0] mem [0:127];
    
    // 读取指令（组合逻辑）
    assign instruction = mem[addr[8:2]];  // 字对齐，忽略低 2 位
    
    // 初始化指令存储器 - 斐波那契数列程序
    // 计算前 10 个斐波那契数并存储到内存
    integer i;
    initial begin
        // 初始化所有指令为 NOP
        for (i = 0; i < 128; i = i + 1) begin
            mem[i] = 32'h00000000;  // NOP (sll $0, $0, 0)
        end
        
        // ===== 6条指令测试程序 =====
        // 测试目标：验证 add, sub, and, or, slt, addi 这6条指令
        // 寄存器使用：
        // $t0 ($8): 测试操作数1 = 5
        // $t1 ($9): 测试操作数2 = 3
        // $t2 ($10): add结果
        // $t3 ($11): sub结果
        // $t4 ($12): and结果
        // $t5 ($13): or结果
        // $t6 ($14): slt结果
        // $t7 ($15): addi结果
        // $s0 ($16): 数据存储基地址 0x100
        
        // 地址 0x00: addi $t0, $0, 7      # $t0 = 7 (测试操作数1)
        mem[0] = 32'h20080007;  // opcode=001000, rs=00000, rt=01000, imm=0000000000000111
        
        // 地址 0x04: addi $t1, $0, 9      # $t1 = 9 (测试操作数2)
        mem[1] = 32'h20090009;  // opcode=001000, rs=00000, rt=01001, imm=0000000000001001
        
        // 地址 0x08: addi $s0, $0, 0x100  # $s0 = 0x100 (数据存储基地址)
        mem[2] = 32'h20100100;  // opcode=001000, rs=00000, rt=10000, imm=0000000100000000
        
        // ===== 测试指令1: add =====
        // 地址 0x0C: add $t2, $t0, $t1    # $t2 = $t0 + $t1 = 5 + 3 = 8
        mem[3] = 32'h01095020;  // opcode=000000, rs=01000, rt=01001, rd=01010, shamt=00000, funct=100000
        
        // 地址 0x10: sw $t2, 0($s0)       # mem[0x100] = $t2 = 8
        mem[4] = 32'hae0a0000;  // opcode=101011, rs=10000, rt=01010, imm=0000000000000000
        
        // ===== 测试指令2: sub =====
        // 地址 0x14: sub $t3, $t0, $t1    # $t3 = $t0 - $t1 = 5 - 3 = 2
        mem[5] = 32'h01095822;  // opcode=000000, rs=01000, rt=01001, rd=01011, shamt=00000, funct=100010
        
        // 地址 0x18: sw $t3, 4($s0)       # mem[0x104] = $t3 = 2
        mem[6] = 32'hae0b0004;  // opcode=101011, rs=10000, rt=01011, imm=0000000000000100
        
        // ===== 测试指令3: and =====
        // 地址 0x1C: and $t4, $t0, $t1    # $t4 = $t0 & $t1 = 5 & 3 = 1
        mem[7] = 32'h01096024;  // opcode=000000, rs=01000, rt=01001, rd=01100, shamt=00000, funct=100100
        
        // 地址 0x20: sw $t4, 8($s0)       # mem[0x108] = $t4 = 1
        mem[8] = 32'hae0c0008;  // opcode=101011, rs=10000, rt=01100, imm=0000000000001000
        
        // ===== 测试指令4: or =====
        // 地址 0x24: or $t5, $t0, $t1     # $t5 = $t0 | $t1 = 5 | 3 = 7
        mem[9] = 32'h01096825;  // opcode=000000, rs=01000, rt=01001, rd=01101, shamt=00000, funct=100101
        
        // 地址 0x28: sw $t5, 12($s0)      # mem[0x10C] = $t5 = 7
        mem[10] = 32'hae0d000c; // opcode=101011, rs=10000, rt=01101, imm=0000000000001100
        
        // ===== 测试指令5: slt =====
        // 地址 0x2C: slt $t6, $t1, $t0    # $t6 = ($t1 < $t0) ? 1 : 0 = (3 < 5) ? 1 : 0 = 1
        mem[11] = 32'h0128702a; // opcode=000000, rs=01001, rt=01000, rd=01110, shamt=00000, funct=101010
        
        // 地址 0x30: sw $t6, 16($s0)      # mem[0x110] = $t6 = 1
        mem[12] = 32'hae0e0010; // opcode=101011, rs=10000, rt=01110, imm=0000000000010000
        
        // ===== 测试指令6: addi =====
        // 地址 0x34: addi $t7, $t0, 10    # $t7 = $t0 + 10 = 5 + 10 = 15
        mem[13] = 32'h210f000a; // opcode=001000, rs=01000, rt=01111, imm=0000000000001010
        
        // 地址 0x38: sw $t7, 20($s0)      # mem[0x114] = $t7 = 15
        mem[14] = 32'hae0f0014; // opcode=101011, rs=10000, rt=01111, imm=0000000000010100
        
        // ===== 验证：使用lw和beq验证结果 =====
        // 地址 0x3C: lw $t8, 0($s0)       # $t8 = mem[0x100] = 8 (验证add结果)
        mem[15] = 32'h8e180000; // opcode=100011, rs=10000, rt=11000, imm=0000000000000000
        
        // 地址 0x40: addi $t9, $0, 8      # $t9 = 8 (期望值)
        mem[16] = 32'h20190008; // opcode=001000, rs=00000, rt=11001, imm=0000000000001000
        
        // 地址 0x44: beq $t8, $t9, 2      # if ($t8 == $t9) 跳转到 END
        mem[17] = 32'h13190002; // opcode=000100, rs=11000, rt=11001, imm=0000000000000010
        
        // 地址 0x48: j 0x50               # 如果验证失败，跳转到错误处理（这里直接跳到结束）
        mem[18] = 32'h08000014; // opcode=000010, addr=00000000000000000000010100
        
        // ===== 程序结束 (END) =====
        // 地址 0x4C: (END标签，无限循环)
        // 地址 0x50: j 0x50               # 无限循环（程序结束）
        mem[20] = 32'h08000014; // opcode=000010, addr=00000000000000000000010100
    end

endmodule
